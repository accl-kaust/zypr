module partial_led_test_v1_0 (
    input clk
);
    
endmodule











































































































































































































































































































































































































