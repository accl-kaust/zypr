
module black_box
(
  input CLK,
  input RST,
  output [7:0] led
);


endmodule
