module thingy (
    input clk,
    output irq
);
    
endmodule







































































































































































































































































































































































































































































































































































































































